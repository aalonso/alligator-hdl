/* wb_gpio.v General pourpuse parallel input/output module
 * Wishbone complaint
 *
 * Copyright (C) 2009 Adrian Alonso Lazcano <aalonso00@gmail.com>
 *
 * This program is free software; you can redistribute it and/or
 * modify it under the terms of the GNU Lesser General Public
 * License as published by the Free Software Foundation; either
 * version 2 of the License, or (at your option) any later version.
 *
 * This program is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU Lesser General Public License for more details.
 *
 * You should have received a copy of the GNU Lesser General Public
 * License along with self library; if not, write to the
 * Free Software Foundation, Inc., 51 Franklin Street, Fifth Floor,
 * Boston, MA 02110-1301, USA.
 *
*/

module wb_gpio (clk_i, rst_i, we_i, stb_i, ack_o, data_i, data_o, irq_o);

	/* TODO add gpio_in gpio_out modules */

endmodule
